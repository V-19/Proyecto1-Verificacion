class stimulus;
  
  rand  logic[31:0] value;//data
  
  rand logic[31:0] value2;//addr
  
  //logic[7:0] bl=($random & 8'h0f)+1;//bl
  
endclass